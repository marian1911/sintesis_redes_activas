** Profile: "SCHEMATIC1-Sim_notch"  [ d:\gd\sintesis de redes activas\sintesis_redes_activas\extra_filtro_notch\filtro_notch-pspicefiles\schematic1\sim_notch.sim ] 

** Creating circuit file "Sim_notch.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\maria\AppData\Roaming\SBP_23.1\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 10 100k
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
