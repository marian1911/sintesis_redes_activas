** Profile: "SCHEMATIC1-Prueba_circ"  [ c:\facultad\materias--4to-2do\sintesis de redes activas\sintesis_redes_activas\tp_balanza\orcad_project\amp_balanza-pspicefiles\schematic1\prueba_circ.sim ] 

** Creating circuit file "Prueba_circ.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\enzog\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1s 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
