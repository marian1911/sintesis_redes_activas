** Profile: "SCHEMATIC1-tp4_montecarlo"  [ D:\GD\Sintesis de redes activas\sintesis_redes_activas\Tp4\tp4_montecarlo-PSpiceFiles\SCHEMATIC1\tp4_montecarlo.sim ] 

** Creating circuit file "tp4_montecarlo.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\maria\AppData\Roaming\SBP_23.1\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 10 1meg
.WCASE AC V([OUT]) YMAX VARY BOTH  HI 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
