** Profile: "SCHEMATIC1-Prueba_circ"  [ d:\gd\sintesis de redes activas\sintesis_redes_activas\tp_balanza\orcad_project\amp_balanza-pspicefiles\schematic1\prueba_circ.sim ] 

** Creating circuit file "Prueba_circ.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\maria\AppData\Roaming\SBP_23.1\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1s 0 
.TEMP 25 125
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
